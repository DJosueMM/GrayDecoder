`timescale 1ns / 1ps

module bin_to_7segmentos_SubModulo( input logic clk,
                                    input logic  [3:0] in,
                                    output logic [6:0] cSeg7);
                                    
    


endmodule
